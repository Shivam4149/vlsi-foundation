module hello;
    initial begin
        $display("VLSI STARTS HERE");
        $finish;
    end
endmodule
