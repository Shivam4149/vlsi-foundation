module hello;
    initial begin
        $display("VLSI GOAT STARTS HERE");
        $finish;
    end
endmodule
